module fc_mac_array #(
   parameter NUM_INPUTS = 48,
   parameter NUM_OUTPUTS = 10,
   parameter DATA_WIDTH = 8,
   parameter ACC_WIDTH = 32
)(
   input clk,
   input rst,
   input valid_in,

   input [DATA_WIDTH*NUM_INPUTS-1:0] data_in_flat,   
   input [DATA_WIDTH*NUM_INPUTS*NUM_OUTPUTS-1:0] weight_flat,

   output reg [ACC_WIDTH*NUM_OUTPUTS-1:0] data_out_flat,   // <-- flat output vector
   output reg finish_sys
);

reg state;
reg [3:0] out_idx;
reg [DATA_WIDTH-1:0] buffer [0:NUM_INPUTS - 1];
reg [DATA_WIDTH - 1:0] weight [0:NUM_INPUTS * NUM_OUTPUTS - 1];

wire [ACC_WIDTH-1:0] calc_out;
reg start_fc;
reg [ACC_WIDTH-1:0] out_reg [0:NUM_OUTPUTS-1];
reg finish_pending;    // <-- added small 1-cycle delay flag

integer i;

always @(posedge clk or posedge rst) begin
   if(rst) begin
      finish_sys <= 0;
      finish_pending <= 0;
      out_idx <= 0;
      state <= 0;
      start_fc <= 0;
      for (i = 0; i < NUM_OUTPUTS; i = i + 1)
         out_reg[i] <= 0;
   end else begin
      if (valid_in)
         start_fc <= 1;

      if(finish_sys == 1)
         finish_sys <= 0;

      if(start_fc == 1) begin
         if(!state) begin
            // unpack 48 inputs from flat vector
            for (i = 0; i < NUM_INPUTS; i = i + 1)
               buffer[i] <= data_in_flat[i*DATA_WIDTH +: DATA_WIDTH];

            // Moved weight unpacking here
            for (i = 0; i < NUM_INPUTS*NUM_OUTPUTS; i = i + 1)
               weight[i] = weight_flat[i*DATA_WIDTH +: DATA_WIDTH];

            state <= 1;
            finish_sys <= 0;
         end else begin
            //out_reg[out_idx] = calc_out;
            out_reg[out_idx] = out_reg[out_idx] + calc_out;
            out_idx <= out_idx + 1'b1;

            if(out_idx == NUM_OUTPUTS) begin
               out_idx <= 0;
               finish_pending <= 1;   // <-- delay finish by 1 cycle
               start_fc <= 0;
               state <= 0;
            end
         end
      end

      // one-cycle delayed flattening
      if (finish_pending) begin
         for (i = 0; i < NUM_OUTPUTS; i = i + 1)
            data_out_flat[i*ACC_WIDTH +: ACC_WIDTH] <= out_reg[i];
         finish_sys <= 1;
         finish_pending <= 0;
      end
   end
end

assign calc_out =
   weight[out_idx * NUM_INPUTS + 0]  * buffer[0]  +
   weight[out_idx * NUM_INPUTS + 1]  * buffer[1]  +
   weight[out_idx * NUM_INPUTS + 2]  * buffer[2]  +
   weight[out_idx * NUM_INPUTS + 3]  * buffer[3]  +
   weight[out_idx * NUM_INPUTS + 4]  * buffer[4]  +
   weight[out_idx * NUM_INPUTS + 5]  * buffer[5]  +
   weight[out_idx * NUM_INPUTS + 6]  * buffer[6]  +
   weight[out_idx * NUM_INPUTS + 7]  * buffer[7]  +
   weight[out_idx * NUM_INPUTS + 8]  * buffer[8]  +
   weight[out_idx * NUM_INPUTS + 9]  * buffer[9]  +
   weight[out_idx * NUM_INPUTS + 10] * buffer[10] +
   weight[out_idx * NUM_INPUTS + 11] * buffer[11] +
   weight[out_idx * NUM_INPUTS + 12] * buffer[12] +
   weight[out_idx * NUM_INPUTS + 13] * buffer[13] +
   weight[out_idx * NUM_INPUTS + 14] * buffer[14] +
   weight[out_idx * NUM_INPUTS + 15] * buffer[15] +
   weight[out_idx * NUM_INPUTS + 16] * buffer[16] +
   weight[out_idx * NUM_INPUTS + 17] * buffer[17] +
   weight[out_idx * NUM_INPUTS + 18] * buffer[18] +
   weight[out_idx * NUM_INPUTS + 19] * buffer[19] +
   weight[out_idx * NUM_INPUTS + 20] * buffer[20] +
   weight[out_idx * NUM_INPUTS + 21] * buffer[21] +
   weight[out_idx * NUM_INPUTS + 22] * buffer[22] +
   weight[out_idx * NUM_INPUTS + 23] * buffer[23] +
   weight[out_idx * NUM_INPUTS + 24] * buffer[24] +
   weight[out_idx * NUM_INPUTS + 25] * buffer[25] +
   weight[out_idx * NUM_INPUTS + 26] * buffer[26] +
   weight[out_idx * NUM_INPUTS + 27] * buffer[27] +
   weight[out_idx * NUM_INPUTS + 28] * buffer[28] +
   weight[out_idx * NUM_INPUTS + 29] * buffer[29] +
   weight[out_idx * NUM_INPUTS + 30] * buffer[30] +
   weight[out_idx * NUM_INPUTS + 31] * buffer[31] +
   weight[out_idx * NUM_INPUTS + 32] * buffer[32] +
   weight[out_idx * NUM_INPUTS + 33] * buffer[33] +
   weight[out_idx * NUM_INPUTS + 34] * buffer[34] +
   weight[out_idx * NUM_INPUTS + 35] * buffer[35] +
   weight[out_idx * NUM_INPUTS + 36] * buffer[36] +
   weight[out_idx * NUM_INPUTS + 37] * buffer[37] +
   weight[out_idx * NUM_INPUTS + 38] * buffer[38] +
   weight[out_idx * NUM_INPUTS + 39] * buffer[39] +
   weight[out_idx * NUM_INPUTS + 40] * buffer[40] +
   weight[out_idx * NUM_INPUTS + 41] * buffer[41] +
   weight[out_idx * NUM_INPUTS + 42] * buffer[42] +
   weight[out_idx * NUM_INPUTS + 43] * buffer[43] +
   weight[out_idx * NUM_INPUTS + 44] * buffer[44] +
   weight[out_idx * NUM_INPUTS + 45] * buffer[45] +
   weight[out_idx * NUM_INPUTS + 46] * buffer[46] +
   weight[out_idx * NUM_INPUTS + 47] * buffer[47];

endmodule
